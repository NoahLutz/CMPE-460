** Profile: "SCHEMATIC1-Csweep"  [ D:\CMPE-460\LABS\Lab7\Lab7-PSpiceFiles\SCHEMATIC1\Csweep.sim ] 

** Creating circuit file "Csweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\cnl9674\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10 1 1e6
.STEP PARAM cap LIST 100e-12 1e-9 10e-9 100e-9 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
